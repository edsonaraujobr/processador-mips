library verilog;
use verilog.vl_types.all;
entity MIPS_VHDL_vlg_vec_tst is
end MIPS_VHDL_vlg_vec_tst;
